-- spi-entity periphiral
-- implements the spi slave
-- 	- handles the miso, mosi
--		- full-duplex => each sck read mosi and write miso

entity spi_entity is 
end entity;

architecture spi_rtl of spi_entity is
begin
end architecture;
