-- fifo-buffer entity
-- implement the fifo buffer handling
-- fifo buffer should reusable for the spi and usb
-- it shouldnt be specifically prepared for either but
-- rather be compatibile with both designs


entity fifo_buffer is
end entity;

architecture fifo_buffer_rtl of fifo_buffer is
begin
end architecture;
