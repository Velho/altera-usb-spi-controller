-- usb-host entity
-- implements the usb host state machine for the ISP1362

entity usb_isp1362_host is
end entity;

architecture rtl_isp1362 of usb_isp1362_host is
begin
end architecture;