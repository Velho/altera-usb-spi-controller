-- top-level vhdl

entity usb_spi_controller is
end entity;

architecture rtl of usb_spi_controller is
begin
end architecture;
